// SoC.v

// Generated using ACDS version 13.1 162 at 2024.04.03.16:26:07

`timescale 1 ps / 1 ps
module SoC (
		input  wire        clk_clk,                            //                         clk.clk
		input  wire        reset_reset_n,                      //                       reset.reset_n
		output wire [2:0]  led_out_external_connection_export, // led_out_external_connection.export
		output wire        pll_c2_clk,                         //                      pll_c2.clk
		output wire [12:0] sdram_controller_wire_addr,         //       sdram_controller_wire.addr
		output wire [1:0]  sdram_controller_wire_ba,           //                            .ba
		output wire        sdram_controller_wire_cas_n,        //                            .cas_n
		output wire        sdram_controller_wire_cke,          //                            .cke
		output wire        sdram_controller_wire_cs_n,         //                            .cs_n
		inout  wire [31:0] sdram_controller_wire_dq,           //                            .dq
		output wire [3:0]  sdram_controller_wire_dqm,          //                            .dqm
		output wire        sdram_controller_wire_ras_n,        //                            .ras_n
		output wire        sdram_controller_wire_we_n          //                            .we_n
	);

	wire         pll_c0_clk;                                                // PLL:c0 -> [CPU:clk, LED_OUT:clk, SDRAM_Controller:clk, clock_crossing_bridge:s0_clk, irq_mapper:clk, irq_synchronizer:sender_clk, jtag_uart:clk, mm_interconnect_1:PLL_c0_clk, rst_controller_001:clk]
	wire         pll_c1_clk;                                                // PLL:c1 -> [SYSID:clock, clock_crossing_bridge:m0_clk, irq_synchronizer:receiver_clk, mm_interconnect_0:PLL_c1_clk, rst_controller_002:clk, timer:clk]
	wire   [0:0] clock_crossing_bridge_m0_burstcount;                       // clock_crossing_bridge:m0_burstcount -> mm_interconnect_0:clock_crossing_bridge_m0_burstcount
	wire         clock_crossing_bridge_m0_waitrequest;                      // mm_interconnect_0:clock_crossing_bridge_m0_waitrequest -> clock_crossing_bridge:m0_waitrequest
	wire   [9:0] clock_crossing_bridge_m0_address;                          // clock_crossing_bridge:m0_address -> mm_interconnect_0:clock_crossing_bridge_m0_address
	wire  [31:0] clock_crossing_bridge_m0_writedata;                        // clock_crossing_bridge:m0_writedata -> mm_interconnect_0:clock_crossing_bridge_m0_writedata
	wire         clock_crossing_bridge_m0_write;                            // clock_crossing_bridge:m0_write -> mm_interconnect_0:clock_crossing_bridge_m0_write
	wire         clock_crossing_bridge_m0_read;                             // clock_crossing_bridge:m0_read -> mm_interconnect_0:clock_crossing_bridge_m0_read
	wire  [31:0] clock_crossing_bridge_m0_readdata;                         // mm_interconnect_0:clock_crossing_bridge_m0_readdata -> clock_crossing_bridge:m0_readdata
	wire         clock_crossing_bridge_m0_debugaccess;                      // clock_crossing_bridge:m0_debugaccess -> mm_interconnect_0:clock_crossing_bridge_m0_debugaccess
	wire   [3:0] clock_crossing_bridge_m0_byteenable;                       // clock_crossing_bridge:m0_byteenable -> mm_interconnect_0:clock_crossing_bridge_m0_byteenable
	wire         clock_crossing_bridge_m0_readdatavalid;                    // mm_interconnect_0:clock_crossing_bridge_m0_readdatavalid -> clock_crossing_bridge:m0_readdatavalid
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:SYSID_control_slave_address -> SYSID:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // SYSID:readdata -> mm_interconnect_0:SYSID_control_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire         mm_interconnect_1_clock_crossing_bridge_s0_waitrequest;    // clock_crossing_bridge:s0_waitrequest -> mm_interconnect_1:clock_crossing_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_1_clock_crossing_bridge_s0_burstcount;     // mm_interconnect_1:clock_crossing_bridge_s0_burstcount -> clock_crossing_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_1_clock_crossing_bridge_s0_writedata;      // mm_interconnect_1:clock_crossing_bridge_s0_writedata -> clock_crossing_bridge:s0_writedata
	wire   [9:0] mm_interconnect_1_clock_crossing_bridge_s0_address;        // mm_interconnect_1:clock_crossing_bridge_s0_address -> clock_crossing_bridge:s0_address
	wire         mm_interconnect_1_clock_crossing_bridge_s0_write;          // mm_interconnect_1:clock_crossing_bridge_s0_write -> clock_crossing_bridge:s0_write
	wire         mm_interconnect_1_clock_crossing_bridge_s0_read;           // mm_interconnect_1:clock_crossing_bridge_s0_read -> clock_crossing_bridge:s0_read
	wire  [31:0] mm_interconnect_1_clock_crossing_bridge_s0_readdata;       // clock_crossing_bridge:s0_readdata -> mm_interconnect_1:clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_1_clock_crossing_bridge_s0_debugaccess;    // mm_interconnect_1:clock_crossing_bridge_s0_debugaccess -> clock_crossing_bridge:s0_debugaccess
	wire         mm_interconnect_1_clock_crossing_bridge_s0_readdatavalid;  // clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_1:clock_crossing_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_clock_crossing_bridge_s0_byteenable;     // mm_interconnect_1:clock_crossing_bridge_s0_byteenable -> clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_1_sdram_controller_s1_waitrequest;         // SDRAM_Controller:za_waitrequest -> mm_interconnect_1:SDRAM_Controller_s1_waitrequest
	wire  [31:0] mm_interconnect_1_sdram_controller_s1_writedata;           // mm_interconnect_1:SDRAM_Controller_s1_writedata -> SDRAM_Controller:az_data
	wire  [24:0] mm_interconnect_1_sdram_controller_s1_address;             // mm_interconnect_1:SDRAM_Controller_s1_address -> SDRAM_Controller:az_addr
	wire         mm_interconnect_1_sdram_controller_s1_chipselect;          // mm_interconnect_1:SDRAM_Controller_s1_chipselect -> SDRAM_Controller:az_cs
	wire         mm_interconnect_1_sdram_controller_s1_write;               // mm_interconnect_1:SDRAM_Controller_s1_write -> SDRAM_Controller:az_wr_n
	wire         mm_interconnect_1_sdram_controller_s1_read;                // mm_interconnect_1:SDRAM_Controller_s1_read -> SDRAM_Controller:az_rd_n
	wire  [31:0] mm_interconnect_1_sdram_controller_s1_readdata;            // SDRAM_Controller:za_data -> mm_interconnect_1:SDRAM_Controller_s1_readdata
	wire         mm_interconnect_1_sdram_controller_s1_readdatavalid;       // SDRAM_Controller:za_valid -> mm_interconnect_1:SDRAM_Controller_s1_readdatavalid
	wire   [3:0] mm_interconnect_1_sdram_controller_s1_byteenable;          // mm_interconnect_1:SDRAM_Controller_s1_byteenable -> SDRAM_Controller:az_be_n
	wire  [31:0] mm_interconnect_1_led_out_s1_writedata;                    // mm_interconnect_1:LED_OUT_s1_writedata -> LED_OUT:writedata
	wire   [1:0] mm_interconnect_1_led_out_s1_address;                      // mm_interconnect_1:LED_OUT_s1_address -> LED_OUT:address
	wire         mm_interconnect_1_led_out_s1_chipselect;                   // mm_interconnect_1:LED_OUT_s1_chipselect -> LED_OUT:chipselect
	wire         mm_interconnect_1_led_out_s1_write;                        // mm_interconnect_1:LED_OUT_s1_write -> LED_OUT:write_n
	wire  [31:0] mm_interconnect_1_led_out_s1_readdata;                     // LED_OUT:readdata -> mm_interconnect_1:LED_OUT_s1_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_1:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                 // CPU:d_writedata -> mm_interconnect_1:CPU_data_master_writedata
	wire  [27:0] cpu_data_master_address;                                   // CPU:d_address -> mm_interconnect_1:CPU_data_master_address
	wire         cpu_data_master_write;                                     // CPU:d_write -> mm_interconnect_1:CPU_data_master_write
	wire         cpu_data_master_read;                                      // CPU:d_read -> mm_interconnect_1:CPU_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_1:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                               // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_1:CPU_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                // CPU:d_byteenable -> mm_interconnect_1:CPU_data_master_byteenable
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_1_pll_pll_slave_writedata;                 // mm_interconnect_1:PLL_pll_slave_writedata -> PLL:writedata
	wire   [1:0] mm_interconnect_1_pll_pll_slave_address;                   // mm_interconnect_1:PLL_pll_slave_address -> PLL:address
	wire         mm_interconnect_1_pll_pll_slave_write;                     // mm_interconnect_1:PLL_pll_slave_write -> PLL:write
	wire         mm_interconnect_1_pll_pll_slave_read;                      // mm_interconnect_1:PLL_pll_slave_read -> PLL:read
	wire  [31:0] mm_interconnect_1_pll_pll_slave_readdata;                  // PLL:readdata -> mm_interconnect_1:PLL_pll_slave_readdata
	wire         mm_interconnect_1_cpu_jtag_debug_module_waitrequest;       // CPU:jtag_debug_module_waitrequest -> mm_interconnect_1:CPU_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_1_cpu_jtag_debug_module_writedata;         // mm_interconnect_1:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_1_cpu_jtag_debug_module_address;           // mm_interconnect_1:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_1_cpu_jtag_debug_module_write;             // mm_interconnect_1:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire         mm_interconnect_1_cpu_jtag_debug_module_read;              // mm_interconnect_1:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire  [31:0] mm_interconnect_1_cpu_jtag_debug_module_readdata;          // CPU:jtag_debug_module_readdata -> mm_interconnect_1:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_1_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_1:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_1_cpu_jtag_debug_module_byteenable;        // mm_interconnect_1:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_1:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // CPU:i_address -> mm_interconnect_1:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                               // CPU:i_read -> mm_interconnect_1:CPU_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_1:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_1:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> CPU:d_irq
	wire         irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                             // timer:irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [PLL:reset, mm_interconnect_1:PLL_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         cpu_jtag_debug_module_reset_reset;                         // CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [CPU:reset_n, LED_OUT:reset_n, SDRAM_Controller:reset_n, clock_crossing_bridge:s0_reset, irq_mapper:reset, irq_synchronizer:sender_reset, jtag_uart:rst_n, mm_interconnect_1:CPU_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [SYSID:reset_n, clock_crossing_bridge:m0_reset, irq_synchronizer:receiver_reset, mm_interconnect_0:clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, timer:reset_n]

	SoC_PLL pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_1_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_1_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_1_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_1_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_1_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (pll_c1_clk),                                //                    c1.clk
		.c2        (pll_c2_clk),                                //                    c2.clk
		.areset    (),                                          //        areset_conduit.export
		.locked    (),                                          //        locked_conduit.export
		.phasedone ()                                           //     phasedone_conduit.export
	);

	SoC_SDRAM_Controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_1_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_1_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_1_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_1_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_1_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_1_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_1_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_1_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_1_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_wire_addr),                          //  wire.export
		.zs_ba          (sdram_controller_wire_ba),                            //      .export
		.zs_cas_n       (sdram_controller_wire_cas_n),                         //      .export
		.zs_cke         (sdram_controller_wire_cke),                           //      .export
		.zs_cs_n        (sdram_controller_wire_cs_n),                          //      .export
		.zs_dq          (sdram_controller_wire_dq),                            //      .export
		.zs_dqm         (sdram_controller_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_controller_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_controller_wire_we_n)                           //      .export
	);

	SoC_timer timer (
		.clk        (pll_c1_clk),                            //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	SoC_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) clock_crossing_bridge (
		.m0_clk           (pll_c1_clk),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                       // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                               //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_1_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_1_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_1_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_1_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_1_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_1_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_1_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_1_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_1_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_1_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	SoC_SYSID sysid (
		.clock    (pll_c1_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	SoC_CPU cpu (
		.clk                                   (pll_c0_clk),                                          //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_1_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_1_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_1_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_1_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_1_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_1_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_1_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_1_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	SoC_LED_OUT led_out (
		.clk        (pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_out_s1_readdata),   //                    .readdata
		.out_port   (led_out_external_connection_export)       // external_connection.export
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.PLL_c1_clk                                                 (pll_c1_clk),                                     //                                               PLL_c1.clk
		.clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),             // clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.clock_crossing_bridge_m0_address                           (clock_crossing_bridge_m0_address),               //                             clock_crossing_bridge_m0.address
		.clock_crossing_bridge_m0_waitrequest                       (clock_crossing_bridge_m0_waitrequest),           //                                                     .waitrequest
		.clock_crossing_bridge_m0_burstcount                        (clock_crossing_bridge_m0_burstcount),            //                                                     .burstcount
		.clock_crossing_bridge_m0_byteenable                        (clock_crossing_bridge_m0_byteenable),            //                                                     .byteenable
		.clock_crossing_bridge_m0_read                              (clock_crossing_bridge_m0_read),                  //                                                     .read
		.clock_crossing_bridge_m0_readdata                          (clock_crossing_bridge_m0_readdata),              //                                                     .readdata
		.clock_crossing_bridge_m0_readdatavalid                     (clock_crossing_bridge_m0_readdatavalid),         //                                                     .readdatavalid
		.clock_crossing_bridge_m0_write                             (clock_crossing_bridge_m0_write),                 //                                                     .write
		.clock_crossing_bridge_m0_writedata                         (clock_crossing_bridge_m0_writedata),             //                                                     .writedata
		.clock_crossing_bridge_m0_debugaccess                       (clock_crossing_bridge_m0_debugaccess),           //                                                     .debugaccess
		.SYSID_control_slave_address                                (mm_interconnect_0_sysid_control_slave_address),  //                                  SYSID_control_slave.address
		.SYSID_control_slave_readdata                               (mm_interconnect_0_sysid_control_slave_readdata), //                                                     .readdata
		.timer_s1_address                                           (mm_interconnect_0_timer_s1_address),             //                                             timer_s1.address
		.timer_s1_write                                             (mm_interconnect_0_timer_s1_write),               //                                                     .write
		.timer_s1_readdata                                          (mm_interconnect_0_timer_s1_readdata),            //                                                     .readdata
		.timer_s1_writedata                                         (mm_interconnect_0_timer_s1_writedata),           //                                                     .writedata
		.timer_s1_chipselect                                        (mm_interconnect_0_timer_s1_chipselect)           //                                                     .chipselect
	);

	SoC_mm_interconnect_1 mm_interconnect_1 (
		.clock_clk_clk                                         (clk_clk),                                                   //                                       clock_clk.clk
		.PLL_c0_clk                                            (pll_c0_clk),                                                //                                          PLL_c0.clk
		.CPU_reset_n_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),                        //               CPU_reset_n_reset_bridge_in_reset.reset
		.PLL_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // PLL_inclk_interface_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                               (cpu_data_master_address),                                   //                                 CPU_data_master.address
		.CPU_data_master_waitrequest                           (cpu_data_master_waitrequest),                               //                                                .waitrequest
		.CPU_data_master_byteenable                            (cpu_data_master_byteenable),                                //                                                .byteenable
		.CPU_data_master_read                                  (cpu_data_master_read),                                      //                                                .read
		.CPU_data_master_readdata                              (cpu_data_master_readdata),                                  //                                                .readdata
		.CPU_data_master_write                                 (cpu_data_master_write),                                     //                                                .write
		.CPU_data_master_writedata                             (cpu_data_master_writedata),                                 //                                                .writedata
		.CPU_data_master_debugaccess                           (cpu_data_master_debugaccess),                               //                                                .debugaccess
		.CPU_instruction_master_address                        (cpu_instruction_master_address),                            //                          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                    (cpu_instruction_master_waitrequest),                        //                                                .waitrequest
		.CPU_instruction_master_read                           (cpu_instruction_master_read),                               //                                                .read
		.CPU_instruction_master_readdata                       (cpu_instruction_master_readdata),                           //                                                .readdata
		.CPU_instruction_master_readdatavalid                  (cpu_instruction_master_readdatavalid),                      //                                                .readdatavalid
		.clock_crossing_bridge_s0_address                      (mm_interconnect_1_clock_crossing_bridge_s0_address),        //                        clock_crossing_bridge_s0.address
		.clock_crossing_bridge_s0_write                        (mm_interconnect_1_clock_crossing_bridge_s0_write),          //                                                .write
		.clock_crossing_bridge_s0_read                         (mm_interconnect_1_clock_crossing_bridge_s0_read),           //                                                .read
		.clock_crossing_bridge_s0_readdata                     (mm_interconnect_1_clock_crossing_bridge_s0_readdata),       //                                                .readdata
		.clock_crossing_bridge_s0_writedata                    (mm_interconnect_1_clock_crossing_bridge_s0_writedata),      //                                                .writedata
		.clock_crossing_bridge_s0_burstcount                   (mm_interconnect_1_clock_crossing_bridge_s0_burstcount),     //                                                .burstcount
		.clock_crossing_bridge_s0_byteenable                   (mm_interconnect_1_clock_crossing_bridge_s0_byteenable),     //                                                .byteenable
		.clock_crossing_bridge_s0_readdatavalid                (mm_interconnect_1_clock_crossing_bridge_s0_readdatavalid),  //                                                .readdatavalid
		.clock_crossing_bridge_s0_waitrequest                  (mm_interconnect_1_clock_crossing_bridge_s0_waitrequest),    //                                                .waitrequest
		.clock_crossing_bridge_s0_debugaccess                  (mm_interconnect_1_clock_crossing_bridge_s0_debugaccess),    //                                                .debugaccess
		.CPU_jtag_debug_module_address                         (mm_interconnect_1_cpu_jtag_debug_module_address),           //                           CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                           (mm_interconnect_1_cpu_jtag_debug_module_write),             //                                                .write
		.CPU_jtag_debug_module_read                            (mm_interconnect_1_cpu_jtag_debug_module_read),              //                                                .read
		.CPU_jtag_debug_module_readdata                        (mm_interconnect_1_cpu_jtag_debug_module_readdata),          //                                                .readdata
		.CPU_jtag_debug_module_writedata                       (mm_interconnect_1_cpu_jtag_debug_module_writedata),         //                                                .writedata
		.CPU_jtag_debug_module_byteenable                      (mm_interconnect_1_cpu_jtag_debug_module_byteenable),        //                                                .byteenable
		.CPU_jtag_debug_module_waitrequest                     (mm_interconnect_1_cpu_jtag_debug_module_waitrequest),       //                                                .waitrequest
		.CPU_jtag_debug_module_debugaccess                     (mm_interconnect_1_cpu_jtag_debug_module_debugaccess),       //                                                .debugaccess
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                .chipselect
		.LED_OUT_s1_address                                    (mm_interconnect_1_led_out_s1_address),                      //                                      LED_OUT_s1.address
		.LED_OUT_s1_write                                      (mm_interconnect_1_led_out_s1_write),                        //                                                .write
		.LED_OUT_s1_readdata                                   (mm_interconnect_1_led_out_s1_readdata),                     //                                                .readdata
		.LED_OUT_s1_writedata                                  (mm_interconnect_1_led_out_s1_writedata),                    //                                                .writedata
		.LED_OUT_s1_chipselect                                 (mm_interconnect_1_led_out_s1_chipselect),                   //                                                .chipselect
		.PLL_pll_slave_address                                 (mm_interconnect_1_pll_pll_slave_address),                   //                                   PLL_pll_slave.address
		.PLL_pll_slave_write                                   (mm_interconnect_1_pll_pll_slave_write),                     //                                                .write
		.PLL_pll_slave_read                                    (mm_interconnect_1_pll_pll_slave_read),                      //                                                .read
		.PLL_pll_slave_readdata                                (mm_interconnect_1_pll_pll_slave_readdata),                  //                                                .readdata
		.PLL_pll_slave_writedata                               (mm_interconnect_1_pll_pll_slave_writedata),                 //                                                .writedata
		.SDRAM_Controller_s1_address                           (mm_interconnect_1_sdram_controller_s1_address),             //                             SDRAM_Controller_s1.address
		.SDRAM_Controller_s1_write                             (mm_interconnect_1_sdram_controller_s1_write),               //                                                .write
		.SDRAM_Controller_s1_read                              (mm_interconnect_1_sdram_controller_s1_read),                //                                                .read
		.SDRAM_Controller_s1_readdata                          (mm_interconnect_1_sdram_controller_s1_readdata),            //                                                .readdata
		.SDRAM_Controller_s1_writedata                         (mm_interconnect_1_sdram_controller_s1_writedata),           //                                                .writedata
		.SDRAM_Controller_s1_byteenable                        (mm_interconnect_1_sdram_controller_s1_byteenable),          //                                                .byteenable
		.SDRAM_Controller_s1_readdatavalid                     (mm_interconnect_1_sdram_controller_s1_readdatavalid),       //                                                .readdatavalid
		.SDRAM_Controller_s1_waitrequest                       (mm_interconnect_1_sdram_controller_s1_waitrequest),         //                                                .waitrequest
		.SDRAM_Controller_s1_chipselect                        (mm_interconnect_1_sdram_controller_s1_chipselect)           //                                                .chipselect
	);

	SoC_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                    // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req      (),                                  // (terminated)
		.reset_req_in0  (1'b0),                              // (terminated)
		.reset_req_in1  (1'b0),                              // (terminated)
		.reset_in2      (1'b0),                              // (terminated)
		.reset_req_in2  (1'b0),                              // (terminated)
		.reset_in3      (1'b0),                              // (terminated)
		.reset_req_in3  (1'b0),                              // (terminated)
		.reset_in4      (1'b0),                              // (terminated)
		.reset_req_in4  (1'b0),                              // (terminated)
		.reset_in5      (1'b0),                              // (terminated)
		.reset_req_in5  (1'b0),                              // (terminated)
		.reset_in6      (1'b0),                              // (terminated)
		.reset_req_in6  (1'b0),                              // (terminated)
		.reset_in7      (1'b0),                              // (terminated)
		.reset_req_in7  (1'b0),                              // (terminated)
		.reset_in8      (1'b0),                              // (terminated)
		.reset_req_in8  (1'b0),                              // (terminated)
		.reset_in9      (1'b0),                              // (terminated)
		.reset_req_in9  (1'b0),                              // (terminated)
		.reset_in10     (1'b0),                              // (terminated)
		.reset_req_in10 (1'b0),                              // (terminated)
		.reset_in11     (1'b0),                              // (terminated)
		.reset_req_in11 (1'b0),                              // (terminated)
		.reset_in12     (1'b0),                              // (terminated)
		.reset_req_in12 (1'b0),                              // (terminated)
		.reset_in13     (1'b0),                              // (terminated)
		.reset_req_in13 (1'b0),                              // (terminated)
		.reset_in14     (1'b0),                              // (terminated)
		.reset_req_in14 (1'b0),                              // (terminated)
		.reset_in15     (1'b0),                              // (terminated)
		.reset_req_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (pll_c1_clk),                         //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
