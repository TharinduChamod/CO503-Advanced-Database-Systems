// SoC.v

// Generated using ACDS version 13.1 162 at 2024.05.22.12:38:02

`timescale 1 ps / 1 ps
module SoC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] mm_interconnect_0_instruction_memory_1_s1_writedata;         // mm_interconnect_0:instruction_memory_1_s1_writedata -> instruction_memory_1:writedata
	wire  [13:0] mm_interconnect_0_instruction_memory_1_s1_address;           // mm_interconnect_0:instruction_memory_1_s1_address -> instruction_memory_1:address
	wire         mm_interconnect_0_instruction_memory_1_s1_chipselect;        // mm_interconnect_0:instruction_memory_1_s1_chipselect -> instruction_memory_1:chipselect
	wire         mm_interconnect_0_instruction_memory_1_s1_clken;             // mm_interconnect_0:instruction_memory_1_s1_clken -> instruction_memory_1:clken
	wire         mm_interconnect_0_instruction_memory_1_s1_write;             // mm_interconnect_0:instruction_memory_1_s1_write -> instruction_memory_1:write
	wire  [31:0] mm_interconnect_0_instruction_memory_1_s1_readdata;          // instruction_memory_1:readdata -> mm_interconnect_0:instruction_memory_1_s1_readdata
	wire   [3:0] mm_interconnect_0_instruction_memory_1_s1_byteenable;        // mm_interconnect_0:instruction_memory_1_s1_byteenable -> instruction_memory_1:byteenable
	wire         cpu_0_data_master_waitrequest;                               // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                 // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [17:0] cpu_0_data_master_address;                                   // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire         cpu_0_data_master_write;                                     // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire         cpu_0_data_master_read;                                      // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire  [31:0] cpu_0_data_master_readdata;                                  // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                               // cpu_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         mm_interconnect_0_fifo_in_waitrequest;                       // FIFO:avalonmm_write_slave_waitrequest -> mm_interconnect_0:FIFO_in_waitrequest
	wire  [31:0] mm_interconnect_0_fifo_in_writedata;                         // mm_interconnect_0:FIFO_in_writedata -> FIFO:avalonmm_write_slave_writedata
	wire         mm_interconnect_0_fifo_in_write;                             // mm_interconnect_0:FIFO_in_write -> FIFO:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_data_memory_0_s1_writedata;                // mm_interconnect_0:data_memory_0_s1_writedata -> data_memory_0:writedata
	wire  [12:0] mm_interconnect_0_data_memory_0_s1_address;                  // mm_interconnect_0:data_memory_0_s1_address -> data_memory_0:address
	wire         mm_interconnect_0_data_memory_0_s1_chipselect;               // mm_interconnect_0:data_memory_0_s1_chipselect -> data_memory_0:chipselect
	wire         mm_interconnect_0_data_memory_0_s1_clken;                    // mm_interconnect_0:data_memory_0_s1_clken -> data_memory_0:clken
	wire         mm_interconnect_0_data_memory_0_s1_write;                    // mm_interconnect_0:data_memory_0_s1_write -> data_memory_0:write
	wire  [31:0] mm_interconnect_0_data_memory_0_s1_readdata;                 // data_memory_0:readdata -> mm_interconnect_0:data_memory_0_s1_readdata
	wire   [3:0] mm_interconnect_0_data_memory_0_s1_byteenable;               // mm_interconnect_0:data_memory_0_s1_byteenable -> data_memory_0:byteenable
	wire         cpu_1_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	wire  [17:0] cpu_1_instruction_master_address;                            // cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	wire         cpu_1_instruction_master_read;                               // cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	wire  [31:0] cpu_1_instruction_master_readdata;                           // mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	wire         cpu_1_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_fifo_out_waitrequest;                      // FIFO:avalonmm_read_slave_waitrequest -> mm_interconnect_0:FIFO_out_waitrequest
	wire         mm_interconnect_0_fifo_out_read;                             // mm_interconnect_0:FIFO_out_read -> FIFO:avalonmm_read_slave_read
	wire  [31:0] mm_interconnect_0_fifo_out_readdata;                         // FIFO:avalonmm_read_slave_readdata -> mm_interconnect_0:FIFO_out_readdata
	wire  [15:0] mm_interconnect_0_highscale_timer_0_s1_writedata;            // mm_interconnect_0:highscale_timer_0_s1_writedata -> highscale_timer_0:writedata
	wire   [2:0] mm_interconnect_0_highscale_timer_0_s1_address;              // mm_interconnect_0:highscale_timer_0_s1_address -> highscale_timer_0:address
	wire         mm_interconnect_0_highscale_timer_0_s1_chipselect;           // mm_interconnect_0:highscale_timer_0_s1_chipselect -> highscale_timer_0:chipselect
	wire         mm_interconnect_0_highscale_timer_0_s1_write;                // mm_interconnect_0:highscale_timer_0_s1_write -> highscale_timer_0:write_n
	wire  [15:0] mm_interconnect_0_highscale_timer_0_s1_readdata;             // highscale_timer_0:readdata -> mm_interconnect_0:highscale_timer_0_s1_readdata
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest; // jtag_uart_1:av_waitrequest -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_writedata -> jtag_uart_1:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_address -> jtag_uart_1:av_address
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_chipselect -> jtag_uart_1:av_chipselect
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_write -> jtag_uart_1:av_write_n
	wire         mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_read -> jtag_uart_1:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata;    // jtag_uart_1:av_readdata -> mm_interconnect_0:jtag_uart_1_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest;       // cpu_1:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_1_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_1_jtag_debug_module_writedata -> cpu_1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_1_jtag_debug_module_address;           // mm_interconnect_0:cpu_1_jtag_debug_module_address -> cpu_1:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_write;             // mm_interconnect_0:cpu_1_jtag_debug_module_write -> cpu_1:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_read;              // mm_interconnect_0:cpu_1_jtag_debug_module_read -> cpu_1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_1_jtag_debug_module_readdata;          // cpu_1:jtag_debug_module_readdata -> mm_interconnect_0:cpu_1_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_1_jtag_debug_module_debugaccess -> cpu_1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_1_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_1_jtag_debug_module_byteenable -> cpu_1:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_highscale_timer_1_s1_writedata;            // mm_interconnect_0:highscale_timer_1_s1_writedata -> highscale_timer_1:writedata
	wire   [2:0] mm_interconnect_0_highscale_timer_1_s1_address;              // mm_interconnect_0:highscale_timer_1_s1_address -> highscale_timer_1:address
	wire         mm_interconnect_0_highscale_timer_1_s1_chipselect;           // mm_interconnect_0:highscale_timer_1_s1_chipselect -> highscale_timer_1:chipselect
	wire         mm_interconnect_0_highscale_timer_1_s1_write;                // mm_interconnect_0:highscale_timer_1_s1_write -> highscale_timer_1:write_n
	wire  [15:0] mm_interconnect_0_highscale_timer_1_s1_readdata;             // highscale_timer_1:readdata -> mm_interconnect_0:highscale_timer_1_s1_readdata
	wire         cpu_1_data_master_waitrequest;                               // mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	wire  [31:0] cpu_1_data_master_writedata;                                 // cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	wire  [17:0] cpu_1_data_master_address;                                   // cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	wire         cpu_1_data_master_write;                                     // cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	wire         cpu_1_data_master_read;                                      // cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	wire  [31:0] cpu_1_data_master_readdata;                                  // mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	wire         cpu_1_data_master_debugaccess;                               // cpu_1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	wire   [3:0] cpu_1_data_master_byteenable;                                // cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	wire  [31:0] mm_interconnect_0_data_memory_1_s1_writedata;                // mm_interconnect_0:data_memory_1_s1_writedata -> data_memory_1:writedata
	wire  [12:0] mm_interconnect_0_data_memory_1_s1_address;                  // mm_interconnect_0:data_memory_1_s1_address -> data_memory_1:address
	wire         mm_interconnect_0_data_memory_1_s1_chipselect;               // mm_interconnect_0:data_memory_1_s1_chipselect -> data_memory_1:chipselect
	wire         mm_interconnect_0_data_memory_1_s1_clken;                    // mm_interconnect_0:data_memory_1_s1_clken -> data_memory_1:clken
	wire         mm_interconnect_0_data_memory_1_s1_write;                    // mm_interconnect_0:data_memory_1_s1_write -> data_memory_1:write
	wire  [31:0] mm_interconnect_0_data_memory_1_s1_readdata;                 // data_memory_1:readdata -> mm_interconnect_0:data_memory_1_s1_readdata
	wire   [3:0] mm_interconnect_0_data_memory_1_s1_byteenable;               // mm_interconnect_0:data_memory_1_s1_byteenable -> data_memory_1:byteenable
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire  [31:0] mm_interconnect_0_instruction_memory_0_s1_writedata;         // mm_interconnect_0:instruction_memory_0_s1_writedata -> instruction_memory_0:writedata
	wire  [13:0] mm_interconnect_0_instruction_memory_0_s1_address;           // mm_interconnect_0:instruction_memory_0_s1_address -> instruction_memory_0:address
	wire         mm_interconnect_0_instruction_memory_0_s1_chipselect;        // mm_interconnect_0:instruction_memory_0_s1_chipselect -> instruction_memory_0:chipselect
	wire         mm_interconnect_0_instruction_memory_0_s1_clken;             // mm_interconnect_0:instruction_memory_0_s1_clken -> instruction_memory_0:clken
	wire         mm_interconnect_0_instruction_memory_0_s1_write;             // mm_interconnect_0:instruction_memory_0_s1_write -> instruction_memory_0:write
	wire  [31:0] mm_interconnect_0_instruction_memory_0_s1_readdata;          // instruction_memory_0:readdata -> mm_interconnect_0:instruction_memory_0_s1_readdata
	wire   [3:0] mm_interconnect_0_instruction_memory_0_s1_byteenable;        // mm_interconnect_0:instruction_memory_0_s1_byteenable -> instruction_memory_0:byteenable
	wire  [31:0] mm_interconnect_0_fifo_in_csr_writedata;                     // mm_interconnect_0:FIFO_in_csr_writedata -> FIFO:wrclk_control_slave_writedata
	wire   [2:0] mm_interconnect_0_fifo_in_csr_address;                       // mm_interconnect_0:FIFO_in_csr_address -> FIFO:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_in_csr_write;                         // mm_interconnect_0:FIFO_in_csr_write -> FIFO:wrclk_control_slave_write
	wire         mm_interconnect_0_fifo_in_csr_read;                          // mm_interconnect_0:FIFO_in_csr_read -> FIFO:wrclk_control_slave_read
	wire  [31:0] mm_interconnect_0_fifo_in_csr_readdata;                      // FIFO:wrclk_control_slave_readdata -> mm_interconnect_0:FIFO_in_csr_readdata
	wire   [0:0] mm_interconnect_0_system_id_control_slave_address;           // mm_interconnect_0:system_id_control_slave_address -> system_id:address
	wire  [31:0] mm_interconnect_0_system_id_control_slave_readdata;          // system_id:readdata -> mm_interconnect_0:system_id_control_slave_readdata
	wire         cpu_0_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [17:0] cpu_0_instruction_master_address;                            // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                               // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire  [31:0] cpu_0_instruction_master_readdata;                           // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest;       // cpu_0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_0_jtag_debug_module_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_0_jtag_debug_module_address;           // mm_interconnect_0:cpu_0_jtag_debug_module_address -> cpu_0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_write;             // mm_interconnect_0:cpu_0_jtag_debug_module_write -> cpu_0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_read;              // mm_interconnect_0:cpu_0_jtag_debug_module_read -> cpu_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_readdata;          // cpu_0:jtag_debug_module_readdata -> mm_interconnect_0:cpu_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_0_jtag_debug_module_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_0_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_0_jtag_debug_module_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver3_irq;                                    // highscale_timer_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_0_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         irq_mapper_001_receiver0_irq;                                // jtag_uart_1:av_irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                // timer_1:irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver3_irq;                                // highscale_timer_1:irq -> irq_mapper_001:receiver3_irq
	wire  [31:0] cpu_1_d_irq_irq;                                             // irq_mapper_001:sender_irq -> cpu_1:d_irq
	wire         irq_mapper_receiver2_irq;                                    // FIFO:wrclk_control_slave_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu_0:reset_n, data_memory_0:reset, highscale_timer_0:reset_n, instruction_memory_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_0_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu_0:reset_req, data_memory_0:reset_req, instruction_memory_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_0_jtag_debug_module_reset_reset;                         // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [FIFO:reset_n, mm_interconnect_0:FIFO_reset_in_reset_bridge_in_reset_reset, system_id:reset_n]
	wire         cpu_1_jtag_debug_module_reset_reset;                         // cpu_1:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in2, rst_controller_002:reset_in1]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [cpu_1:reset_n, data_memory_1:reset, highscale_timer_1:reset_n, instruction_memory_1:reset, irq_mapper_001:reset, jtag_uart_1:rst_n, mm_interconnect_0:cpu_1_reset_n_reset_bridge_in_reset_reset, rst_translator_001:in_reset, timer_1:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [cpu_1:reset_req, data_memory_1:reset_req, instruction_memory_1:reset_req, rst_translator_001:reset_req_in]

	SoC_cpu_0 cpu_0 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (cpu_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_0_data_master_read),                                //                          .read
		.d_readdata                            (cpu_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_0_data_master_write),                               //                          .write
		.d_writedata                           (cpu_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	SoC_instruction_memory_0 instruction_memory_0 (
		.clk        (clk_clk),                                              //   clk1.clk
		.address    (mm_interconnect_0_instruction_memory_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_instruction_memory_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_instruction_memory_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_instruction_memory_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_instruction_memory_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_instruction_memory_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_instruction_memory_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                    //       .reset_req
	);

	SoC_data_memory_0 data_memory_0 (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_data_memory_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	SoC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	SoC_system_id system_id (
		.clock    (clk_clk),                                            //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_system_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_system_id_control_slave_address)   //              .address
	);

	SoC_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	SoC_cpu_1 cpu_1 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                   //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),                //                          .reset_req
		.d_address                             (cpu_1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_1_data_master_read),                                //                          .read
		.d_readdata                            (cpu_1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_1_data_master_write),                               //                          .write
		.d_writedata                           (cpu_1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_1_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_1_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_1_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	SoC_instruction_memory_1 instruction_memory_1 (
		.clk        (clk_clk),                                              //   clk1.clk
		.address    (mm_interconnect_0_instruction_memory_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_instruction_memory_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_instruction_memory_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_instruction_memory_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_instruction_memory_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_instruction_memory_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_instruction_memory_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)                //       .reset_req
	);

	SoC_data_memory_1 data_memory_1 (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_data_memory_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)         //       .reset_req
	);

	SoC_jtag_uart_0 jtag_uart_1 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver0_irq)                                 //               irq.irq
	);

	SoC_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver1_irq)             //   irq.irq
	);

	SoC_FIFO fifo (
		.wrclock                          (clk_clk),                                 //   clk_in.clk
		.reset_n                          (~rst_controller_001_reset_out_reset),     // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_fifo_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_fifo_in_write),         //         .write
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_fifo_in_waitrequest),   //         .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_out_read),         //         .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address      (mm_interconnect_0_fifo_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_fifo_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_fifo_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_fifo_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_fifo_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver2_irq)                 //   in_irq.irq
	);

	SoC_highscale_timer_0 highscale_timer_0 (
		.clk        (clk_clk),                                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   // reset.reset_n
		.address    (mm_interconnect_0_highscale_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_highscale_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_highscale_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_highscale_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_highscale_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                           //   irq.irq
	);

	SoC_highscale_timer_0 highscale_timer_1 (
		.clk        (clk_clk),                                           //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_highscale_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_highscale_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_highscale_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_highscale_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_highscale_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver3_irq)                       //   irq.irq
	);

	SoC_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                             (clk_clk),                                                     //                           clock_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // cpu_0_reset_n_reset_bridge_in_reset.reset
		.cpu_1_reset_n_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // cpu_1_reset_n_reset_bridge_in_reset.reset
		.FIFO_reset_in_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // FIFO_reset_in_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                 (cpu_0_data_master_address),                                   //                   cpu_0_data_master.address
		.cpu_0_data_master_waitrequest             (cpu_0_data_master_waitrequest),                               //                                    .waitrequest
		.cpu_0_data_master_byteenable              (cpu_0_data_master_byteenable),                                //                                    .byteenable
		.cpu_0_data_master_read                    (cpu_0_data_master_read),                                      //                                    .read
		.cpu_0_data_master_readdata                (cpu_0_data_master_readdata),                                  //                                    .readdata
		.cpu_0_data_master_write                   (cpu_0_data_master_write),                                     //                                    .write
		.cpu_0_data_master_writedata               (cpu_0_data_master_writedata),                                 //                                    .writedata
		.cpu_0_data_master_debugaccess             (cpu_0_data_master_debugaccess),                               //                                    .debugaccess
		.cpu_0_instruction_master_address          (cpu_0_instruction_master_address),                            //            cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest      (cpu_0_instruction_master_waitrequest),                        //                                    .waitrequest
		.cpu_0_instruction_master_read             (cpu_0_instruction_master_read),                               //                                    .read
		.cpu_0_instruction_master_readdata         (cpu_0_instruction_master_readdata),                           //                                    .readdata
		.cpu_0_instruction_master_readdatavalid    (cpu_0_instruction_master_readdatavalid),                      //                                    .readdatavalid
		.cpu_1_data_master_address                 (cpu_1_data_master_address),                                   //                   cpu_1_data_master.address
		.cpu_1_data_master_waitrequest             (cpu_1_data_master_waitrequest),                               //                                    .waitrequest
		.cpu_1_data_master_byteenable              (cpu_1_data_master_byteenable),                                //                                    .byteenable
		.cpu_1_data_master_read                    (cpu_1_data_master_read),                                      //                                    .read
		.cpu_1_data_master_readdata                (cpu_1_data_master_readdata),                                  //                                    .readdata
		.cpu_1_data_master_write                   (cpu_1_data_master_write),                                     //                                    .write
		.cpu_1_data_master_writedata               (cpu_1_data_master_writedata),                                 //                                    .writedata
		.cpu_1_data_master_debugaccess             (cpu_1_data_master_debugaccess),                               //                                    .debugaccess
		.cpu_1_instruction_master_address          (cpu_1_instruction_master_address),                            //            cpu_1_instruction_master.address
		.cpu_1_instruction_master_waitrequest      (cpu_1_instruction_master_waitrequest),                        //                                    .waitrequest
		.cpu_1_instruction_master_read             (cpu_1_instruction_master_read),                               //                                    .read
		.cpu_1_instruction_master_readdata         (cpu_1_instruction_master_readdata),                           //                                    .readdata
		.cpu_1_instruction_master_readdatavalid    (cpu_1_instruction_master_readdatavalid),                      //                                    .readdatavalid
		.cpu_0_jtag_debug_module_address           (mm_interconnect_0_cpu_0_jtag_debug_module_address),           //             cpu_0_jtag_debug_module.address
		.cpu_0_jtag_debug_module_write             (mm_interconnect_0_cpu_0_jtag_debug_module_write),             //                                    .write
		.cpu_0_jtag_debug_module_read              (mm_interconnect_0_cpu_0_jtag_debug_module_read),              //                                    .read
		.cpu_0_jtag_debug_module_readdata          (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),          //                                    .readdata
		.cpu_0_jtag_debug_module_writedata         (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),         //                                    .writedata
		.cpu_0_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),        //                                    .byteenable
		.cpu_0_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest),       //                                    .waitrequest
		.cpu_0_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess),       //                                    .debugaccess
		.cpu_1_jtag_debug_module_address           (mm_interconnect_0_cpu_1_jtag_debug_module_address),           //             cpu_1_jtag_debug_module.address
		.cpu_1_jtag_debug_module_write             (mm_interconnect_0_cpu_1_jtag_debug_module_write),             //                                    .write
		.cpu_1_jtag_debug_module_read              (mm_interconnect_0_cpu_1_jtag_debug_module_read),              //                                    .read
		.cpu_1_jtag_debug_module_readdata          (mm_interconnect_0_cpu_1_jtag_debug_module_readdata),          //                                    .readdata
		.cpu_1_jtag_debug_module_writedata         (mm_interconnect_0_cpu_1_jtag_debug_module_writedata),         //                                    .writedata
		.cpu_1_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_1_jtag_debug_module_byteenable),        //                                    .byteenable
		.cpu_1_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_1_jtag_debug_module_waitrequest),       //                                    .waitrequest
		.cpu_1_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_1_jtag_debug_module_debugaccess),       //                                    .debugaccess
		.data_memory_0_s1_address                  (mm_interconnect_0_data_memory_0_s1_address),                  //                    data_memory_0_s1.address
		.data_memory_0_s1_write                    (mm_interconnect_0_data_memory_0_s1_write),                    //                                    .write
		.data_memory_0_s1_readdata                 (mm_interconnect_0_data_memory_0_s1_readdata),                 //                                    .readdata
		.data_memory_0_s1_writedata                (mm_interconnect_0_data_memory_0_s1_writedata),                //                                    .writedata
		.data_memory_0_s1_byteenable               (mm_interconnect_0_data_memory_0_s1_byteenable),               //                                    .byteenable
		.data_memory_0_s1_chipselect               (mm_interconnect_0_data_memory_0_s1_chipselect),               //                                    .chipselect
		.data_memory_0_s1_clken                    (mm_interconnect_0_data_memory_0_s1_clken),                    //                                    .clken
		.data_memory_1_s1_address                  (mm_interconnect_0_data_memory_1_s1_address),                  //                    data_memory_1_s1.address
		.data_memory_1_s1_write                    (mm_interconnect_0_data_memory_1_s1_write),                    //                                    .write
		.data_memory_1_s1_readdata                 (mm_interconnect_0_data_memory_1_s1_readdata),                 //                                    .readdata
		.data_memory_1_s1_writedata                (mm_interconnect_0_data_memory_1_s1_writedata),                //                                    .writedata
		.data_memory_1_s1_byteenable               (mm_interconnect_0_data_memory_1_s1_byteenable),               //                                    .byteenable
		.data_memory_1_s1_chipselect               (mm_interconnect_0_data_memory_1_s1_chipselect),               //                                    .chipselect
		.data_memory_1_s1_clken                    (mm_interconnect_0_data_memory_1_s1_clken),                    //                                    .clken
		.FIFO_in_write                             (mm_interconnect_0_fifo_in_write),                             //                             FIFO_in.write
		.FIFO_in_writedata                         (mm_interconnect_0_fifo_in_writedata),                         //                                    .writedata
		.FIFO_in_waitrequest                       (mm_interconnect_0_fifo_in_waitrequest),                       //                                    .waitrequest
		.FIFO_in_csr_address                       (mm_interconnect_0_fifo_in_csr_address),                       //                         FIFO_in_csr.address
		.FIFO_in_csr_write                         (mm_interconnect_0_fifo_in_csr_write),                         //                                    .write
		.FIFO_in_csr_read                          (mm_interconnect_0_fifo_in_csr_read),                          //                                    .read
		.FIFO_in_csr_readdata                      (mm_interconnect_0_fifo_in_csr_readdata),                      //                                    .readdata
		.FIFO_in_csr_writedata                     (mm_interconnect_0_fifo_in_csr_writedata),                     //                                    .writedata
		.FIFO_out_read                             (mm_interconnect_0_fifo_out_read),                             //                            FIFO_out.read
		.FIFO_out_readdata                         (mm_interconnect_0_fifo_out_readdata),                         //                                    .readdata
		.FIFO_out_waitrequest                      (mm_interconnect_0_fifo_out_waitrequest),                      //                                    .waitrequest
		.highscale_timer_0_s1_address              (mm_interconnect_0_highscale_timer_0_s1_address),              //                highscale_timer_0_s1.address
		.highscale_timer_0_s1_write                (mm_interconnect_0_highscale_timer_0_s1_write),                //                                    .write
		.highscale_timer_0_s1_readdata             (mm_interconnect_0_highscale_timer_0_s1_readdata),             //                                    .readdata
		.highscale_timer_0_s1_writedata            (mm_interconnect_0_highscale_timer_0_s1_writedata),            //                                    .writedata
		.highscale_timer_0_s1_chipselect           (mm_interconnect_0_highscale_timer_0_s1_chipselect),           //                                    .chipselect
		.highscale_timer_1_s1_address              (mm_interconnect_0_highscale_timer_1_s1_address),              //                highscale_timer_1_s1.address
		.highscale_timer_1_s1_write                (mm_interconnect_0_highscale_timer_1_s1_write),                //                                    .write
		.highscale_timer_1_s1_readdata             (mm_interconnect_0_highscale_timer_1_s1_readdata),             //                                    .readdata
		.highscale_timer_1_s1_writedata            (mm_interconnect_0_highscale_timer_1_s1_writedata),            //                                    .writedata
		.highscale_timer_1_s1_chipselect           (mm_interconnect_0_highscale_timer_1_s1_chipselect),           //                                    .chipselect
		.instruction_memory_0_s1_address           (mm_interconnect_0_instruction_memory_0_s1_address),           //             instruction_memory_0_s1.address
		.instruction_memory_0_s1_write             (mm_interconnect_0_instruction_memory_0_s1_write),             //                                    .write
		.instruction_memory_0_s1_readdata          (mm_interconnect_0_instruction_memory_0_s1_readdata),          //                                    .readdata
		.instruction_memory_0_s1_writedata         (mm_interconnect_0_instruction_memory_0_s1_writedata),         //                                    .writedata
		.instruction_memory_0_s1_byteenable        (mm_interconnect_0_instruction_memory_0_s1_byteenable),        //                                    .byteenable
		.instruction_memory_0_s1_chipselect        (mm_interconnect_0_instruction_memory_0_s1_chipselect),        //                                    .chipselect
		.instruction_memory_0_s1_clken             (mm_interconnect_0_instruction_memory_0_s1_clken),             //                                    .clken
		.instruction_memory_1_s1_address           (mm_interconnect_0_instruction_memory_1_s1_address),           //             instruction_memory_1_s1.address
		.instruction_memory_1_s1_write             (mm_interconnect_0_instruction_memory_1_s1_write),             //                                    .write
		.instruction_memory_1_s1_readdata          (mm_interconnect_0_instruction_memory_1_s1_readdata),          //                                    .readdata
		.instruction_memory_1_s1_writedata         (mm_interconnect_0_instruction_memory_1_s1_writedata),         //                                    .writedata
		.instruction_memory_1_s1_byteenable        (mm_interconnect_0_instruction_memory_1_s1_byteenable),        //                                    .byteenable
		.instruction_memory_1_s1_chipselect        (mm_interconnect_0_instruction_memory_1_s1_chipselect),        //                                    .chipselect
		.instruction_memory_1_s1_clken             (mm_interconnect_0_instruction_memory_1_s1_clken),             //                                    .clken
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.jtag_uart_1_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_address),     //       jtag_uart_1_avalon_jtag_slave.address
		.jtag_uart_1_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_1_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_1_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_1_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_1_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_1_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_1_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.system_id_control_slave_address           (mm_interconnect_0_system_id_control_slave_address),           //             system_id_control_slave.address
		.system_id_control_slave_readdata          (mm_interconnect_0_system_id_control_slave_readdata),          //                                    .readdata
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                        //                          timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                          //                                    .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                       //                                    .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),                      //                                    .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect),                     //                                    .chipselect
		.timer_1_s1_address                        (mm_interconnect_0_timer_1_s1_address),                        //                          timer_1_s1.address
		.timer_1_s1_write                          (mm_interconnect_0_timer_1_s1_write),                          //                                    .write
		.timer_1_s1_readdata                       (mm_interconnect_0_timer_1_s1_readdata),                       //                                    .readdata
		.timer_1_s1_writedata                      (mm_interconnect_0_timer_1_s1_writedata),                      //                                    .writedata
		.timer_1_s1_chipselect                     (mm_interconnect_0_timer_1_s1_chipselect)                      //                                    .chipselect
	);

	SoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	SoC_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_1_d_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (cpu_1_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_1_jtag_debug_module_reset_reset),    // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
